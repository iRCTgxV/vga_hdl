// clock_108Mhz.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module clock_108Mhz (
		input  wire  clk_in_clk,         //         clk_in.clk
		output wire  clk_out_108mhz_clk, // clk_out_108mhz.clk
		input  wire  rst_reset           //            rst.reset
	);

	clock_108Mhz_pll_0 pll_0 (
		.refclk   (clk_in_clk),         //  refclk.clk
		.rst      (rst_reset),          //   reset.reset
		.outclk_0 (clk_out_108mhz_clk), // outclk0.clk
		.locked   ()                    // (terminated)
	);

endmodule
