
module clock_108Mhz (
	clk_in_clk,
	rst_reset,
	clk_out_108mhz_clk);	

	input		clk_in_clk;
	input		rst_reset;
	output		clk_out_108mhz_clk;
endmodule
